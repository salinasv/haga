
--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   19:43:17 09/30/2008
-- Design Name:   order_perm
-- Module Name:   /home/salinasv/George/George/1Ise/Tesis/Xilinx/TSP_SEP_27/tb_order_perm.vhd
-- Project Name:  TSP_SEP_27
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: order_perm
--
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends 
-- that these types always be used for the top-level I/O of a design in order 
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_arith.ALL;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.ALL;

ENTITY tb_order_perm_vhd IS
END tb_order_perm_vhd;

ARCHITECTURE behavior OF tb_order_perm_vhd IS 

	-- Component Declaration for the Unit Under Test (UUT)
	COMPONENT order_perm
	generic (
		DATA_WIDTH	: integer;	-- natural register size
		M_LOG2		: integer		-- log2(m)
	);
	PORT(
		clk : IN std_logic;
		Dat_in : IN std_logic_vector(7 downto 0);
		reset : IN std_logic;
		datram : OUT std_logic_vector(7 downto 0);
		addr : OUT std_logic_vector(7 downto 0);
		WE : OUT std_logic;
		Done : OUT std_logic
		);
	END COMPONENT;

	--Inputs
	SIGNAL clk :  std_logic := '0';
	SIGNAL reset :  std_logic := '1';
	SIGNAL Dat_in :  std_logic_vector(7 downto 0) := (others=>'0');

	--Outputs
	SIGNAL Datram : std_logic_vector(7 downto 0) := (others => '0');
	SIGNAL addr :  std_logic_vector(7 downto 0) := (others => '0');
	SIGNAL WE :  std_logic := '0';
	SIGNAL Done :  std_logic := '0';

	constant clk_T : time := 3 ns;
	--signal iter : std_logic_vector(8-1 downto 0) := 254; --(others => '1');
	signal iter : integer range 0 to 256 := 255; --(others => '1');
	--constant LAST : std_logic_vector(8-1 downto 0) := (others => '1');
	constant LAST : integer := 256;
	signal perm_data : integer := 0;
	
	type perm_ram_type is array (0 to (10*(2**8))-1) of integer;
	signal ram_out : perm_ram_type := (others => 0);

	constant perm_rom : perm_ram_type :=
	(
175, 31, 12, 3, 185, 54, 183, 72, 71, 122, 0, 148, 187, 74, 68, 203, 151, 219, 49, 66, 179, 204, 26, 125, 177, 56, 193, 190, 225, 139, 7, 92, 2, 152, 221, 166, 118, 255, 206, 19, 23, 76, 103, 111, 42, 254, 250, 28, 140, 209, 17, 130, 145, 13, 6, 117, 79, 136, 11, 253, 32, 75, 67, 252, 157, 27, 218, 233, 25, 138, 61, 142, 189, 126, 172, 160, 63, 153, 199, 96, 22, 93, 176, 147, 50, 195, 107, 197, 213, 38, 243, 18, 178, 37, 123, 244, 214, 114, 205, 24, 239, 94, 124, 36, 246, 101, 90, 201, 109, 222, 10, 245, 80, 108, 89, 59, 112, 182, 53, 110, 236, 150, 235, 141, 128, 105, 60, 224, 154, 85, 165, 161, 216, 192, 86, 116, 228, 35, 95, 220, 100, 82, 196, 81, 45, 21, 15, 242, 158, 70, 170, 226, 69, 62, 88, 29, 171, 230, 64, 188, 99, 20, 84, 47, 91, 33, 57, 102, 247, 98, 4, 237, 234, 43, 14, 249, 200, 30, 223, 46, 78, 40, 146, 251, 34, 97, 65, 132, 106, 238, 44, 211, 144, 184, 163, 55, 180, 217, 210, 1, 202, 191, 120, 51, 48, 162, 215, 212, 77, 119, 129, 127, 159, 229, 169, 121, 58, 39, 227, 83, 241, 231, 248, 16, 186, 41, 52, 173, 207, 8, 194, 133, 137, 134, 174, 156, 198, 104, 135, 131, 9, 164, 149, 87, 181, 240, 155, 113, 5, 167, 208, 232, 73, 115, 168, 143, 
136, 167, 141, 146, 64, 37, 99, 202, 219, 16, 47, 28, 254, 126, 78, 83, 48, 197, 220, 86, 182, 253, 90, 169, 30, 31, 104, 135, 38, 212, 149, 108, 139, 200, 155, 238, 116, 7, 244, 143, 243, 234, 119, 138, 123, 162, 175, 26, 185, 230, 92, 144, 181, 142, 152, 228, 67, 125, 160, 4, 188, 69, 46, 65, 158, 115, 163, 58, 124, 170, 164, 221, 41, 20, 168, 0, 109, 61, 29, 232, 229, 209, 62, 79, 255, 117, 60, 50, 18, 172, 241, 194, 248, 27, 195, 184, 44, 98, 77, 251, 52, 76, 10, 89, 45, 129, 236, 190, 25, 121, 39, 51, 193, 53, 246, 199, 215, 247, 140, 111, 208, 156, 56, 35, 14, 80, 187, 17, 102, 5, 75, 174, 63, 94, 68, 96, 206, 97, 43, 36, 42, 176, 23, 82, 252, 165, 191, 1, 8, 240, 214, 203, 249, 250, 137, 13, 171, 132, 154, 210, 201, 106, 222, 107, 178, 93, 211, 186, 21, 2, 22, 110, 231, 150, 196, 81, 213, 32, 103, 40, 19, 216, 59, 54, 173, 189, 33, 122, 177, 24, 218, 180, 71, 161, 223, 217, 245, 72, 148, 131, 70, 198, 118, 55, 145, 114, 57, 113, 147, 235, 66, 204, 239, 101, 73, 205, 151, 128, 85, 105, 127, 159, 179, 134, 91, 224, 34, 227, 3, 12, 11, 9, 120, 242, 15, 153, 207, 225, 183, 95, 49, 133, 157, 112, 6, 84, 100, 233, 237, 88, 166, 130, 74, 87, 226, 192, 
17, 67, 119, 124, 34, 111, 135, 197, 182, 59, 148, 23, 235, 7, 164, 227, 83, 122, 156, 74, 97, 31, 73, 189, 61, 239, 230, 171, 68, 199, 99, 221, 58, 47, 123, 242, 56, 81, 180, 66, 126, 225, 42, 193, 9, 79, 53, 161, 22, 8, 48, 228, 24, 179, 167, 237, 162, 29, 245, 254, 76, 32, 105, 240, 248, 195, 213, 13, 232, 198, 142, 175, 191, 154, 192, 155, 121, 140, 146, 214, 118, 4, 86, 38, 40, 41, 130, 204, 80, 166, 209, 127, 117, 95, 168, 12, 77, 158, 149, 72, 33, 51, 102, 94, 203, 2, 27, 110, 176, 30, 129, 201, 112, 205, 114, 251, 16, 52, 177, 141, 224, 220, 55, 64, 188, 116, 93, 19, 194, 54, 160, 196, 253, 133, 91, 87, 115, 165, 138, 241, 206, 139, 212, 137, 200, 49, 247, 25, 229, 222, 120, 5, 36, 147, 109, 134, 249, 208, 226, 0, 92, 252, 202, 184, 152, 217, 45, 173, 50, 132, 101, 26, 37, 143, 187, 71, 10, 75, 159, 210, 234, 46, 244, 246, 35, 113, 69, 96, 172, 89, 231, 128, 170, 43, 211, 144, 207, 233, 181, 103, 153, 39, 20, 82, 62, 21, 84, 216, 151, 6, 106, 183, 219, 157, 14, 90, 100, 11, 57, 178, 190, 131, 15, 65, 243, 60, 1, 186, 185, 88, 223, 136, 236, 145, 215, 3, 98, 255, 18, 63, 238, 150, 85, 169, 107, 78, 163, 108, 70, 174, 104, 250, 28, 44, 125, 218, 
91, 72, 210, 199, 64, 84, 81, 129, 105, 207, 240, 183, 153, 204, 163, 78, 60, 171, 137, 82, 57, 77, 146, 231, 71, 132, 203, 190, 250, 120, 25, 80, 1, 66, 172, 10, 18, 43, 131, 202, 255, 140, 119, 242, 104, 112, 116, 4, 94, 110, 232, 73, 200, 127, 30, 55, 196, 253, 123, 228, 97, 181, 90, 26, 35, 68, 93, 67, 151, 59, 152, 122, 184, 194, 16, 221, 39, 54, 219, 212, 34, 98, 206, 238, 154, 50, 213, 89, 128, 99, 107, 176, 244, 41, 13, 75, 6, 177, 189, 86, 118, 85, 126, 79, 133, 111, 157, 158, 53, 51, 248, 252, 178, 168, 226, 162, 245, 205, 95, 103, 96, 167, 254, 37, 201, 138, 243, 193, 88, 65, 42, 32, 145, 24, 7, 147, 2, 45, 230, 247, 70, 121, 237, 44, 38, 100, 87, 208, 28, 141, 20, 179, 155, 27, 29, 209, 239, 218, 11, 0, 175, 160, 108, 76, 69, 63, 9, 220, 48, 161, 249, 229, 125, 15, 36, 62, 61, 143, 215, 149, 92, 182, 166, 170, 165, 33, 191, 139, 142, 114, 197, 74, 46, 159, 134, 222, 124, 173, 117, 21, 235, 187, 102, 109, 251, 49, 185, 211, 188, 234, 150, 17, 241, 113, 246, 223, 135, 136, 192, 115, 144, 52, 47, 174, 40, 217, 14, 56, 164, 169, 214, 180, 236, 101, 156, 148, 198, 225, 227, 23, 22, 216, 195, 3, 19, 233, 106, 5, 12, 83, 130, 186, 58, 31, 8, 224, 
34, 6, 252, 200, 191, 74, 15, 97, 230, 138, 192, 165, 124, 35, 3, 169, 50, 30, 0, 142, 239, 103, 21, 210, 137, 32, 216, 17, 101, 66, 79, 52, 98, 198, 197, 117, 232, 246, 149, 193, 180, 61, 109, 217, 160, 23, 70, 144, 212, 33, 159, 199, 238, 167, 206, 154, 128, 9, 214, 223, 46, 106, 56, 83, 119, 158, 196, 107, 45, 94, 65, 255, 162, 81, 249, 133, 110, 122, 71, 113, 233, 175, 155, 39, 135, 76, 222, 38, 136, 134, 25, 152, 211, 208, 77, 96, 182, 99, 14, 40, 242, 100, 139, 118, 53, 41, 80, 75, 181, 150, 185, 115, 36, 204, 69, 245, 114, 49, 171, 178, 163, 7, 228, 243, 221, 18, 241, 78, 190, 179, 195, 125, 58, 201, 102, 22, 253, 130, 166, 64, 95, 12, 188, 224, 73, 244, 189, 10, 247, 157, 131, 161, 108, 240, 59, 60, 4, 132, 254, 29, 126, 236, 20, 164, 176, 235, 231, 62, 54, 120, 213, 90, 111, 116, 156, 148, 93, 57, 177, 27, 218, 92, 207, 47, 72, 26, 82, 234, 37, 194, 143, 121, 172, 87, 5, 16, 205, 225, 209, 1, 112, 55, 8, 251, 44, 147, 19, 11, 28, 203, 220, 31, 145, 86, 237, 202, 183, 229, 24, 227, 91, 184, 226, 13, 123, 48, 104, 43, 168, 219, 42, 146, 173, 51, 186, 84, 170, 88, 63, 250, 2, 67, 174, 85, 129, 215, 68, 140, 151, 141, 153, 187, 248, 127, 89, 105, 
215, 67, 95, 26, 81, 29, 141, 74, 65, 129, 136, 166, 133, 1, 9, 177, 125, 93, 62, 55, 36, 172, 240, 207, 139, 42, 92, 11, 2, 204, 233, 244, 31, 247, 185, 69, 59, 84, 76, 28, 21, 181, 24, 78, 239, 46, 254, 53, 248, 63, 173, 205, 249, 255, 243, 56, 217, 161, 50, 12, 140, 228, 188, 117, 150, 75, 175, 100, 196, 187, 182, 198, 10, 54, 49, 218, 223, 109, 145, 73, 88, 77, 51, 90, 94, 82, 45, 58, 227, 87, 192, 153, 199, 203, 115, 167, 38, 124, 253, 246, 0, 220, 168, 70, 206, 202, 211, 22, 245, 128, 43, 83, 34, 18, 221, 230, 214, 226, 212, 114, 122, 222, 123, 130, 200, 107, 33, 183, 41, 86, 208, 252, 157, 231, 66, 156, 169, 229, 195, 176, 68, 170, 178, 152, 190, 60, 91, 209, 52, 16, 13, 180, 47, 146, 158, 64, 151, 154, 44, 232, 103, 101, 225, 142, 164, 113, 219, 80, 108, 57, 30, 201, 235, 241, 48, 104, 112, 20, 99, 165, 102, 162, 121, 98, 111, 191, 186, 236, 7, 79, 14, 3, 189, 143, 23, 179, 19, 138, 27, 106, 61, 126, 4, 250, 120, 118, 159, 174, 193, 37, 97, 194, 210, 216, 184, 71, 144, 17, 85, 213, 116, 32, 148, 15, 96, 35, 132, 238, 8, 39, 72, 171, 251, 197, 40, 25, 149, 160, 224, 242, 137, 163, 6, 105, 89, 131, 127, 135, 155, 237, 234, 134, 119, 147, 110, 5, 
219, 187, 122, 104, 6, 4, 5, 93, 67, 182, 18, 51, 246, 108, 158, 74, 139, 59, 10, 253, 56, 201, 192, 135, 117, 211, 179, 105, 22, 99, 109, 183, 198, 238, 239, 29, 237, 7, 255, 184, 140, 62, 119, 230, 98, 142, 132, 254, 202, 17, 90, 63, 45, 20, 159, 163, 188, 40, 229, 245, 64, 150, 148, 76, 164, 111, 26, 86, 75, 213, 249, 180, 177, 251, 137, 240, 80, 170, 121, 118, 126, 168, 220, 39, 200, 243, 120, 44, 94, 2, 236, 156, 31, 134, 78, 131, 216, 167, 214, 46, 125, 16, 169, 161, 145, 146, 244, 82, 12, 133, 89, 103, 54, 8, 107, 42, 13, 155, 223, 50, 233, 24, 60, 33, 199, 181, 87, 21, 43, 124, 49, 191, 221, 11, 115, 1, 152, 61, 97, 27, 196, 79, 100, 0, 32, 250, 130, 19, 189, 57, 83, 95, 203, 197, 208, 174, 194, 106, 235, 41, 160, 96, 154, 30, 9, 129, 173, 228, 232, 36, 69, 35, 205, 153, 176, 186, 209, 127, 149, 25, 114, 88, 207, 68, 110, 225, 38, 34, 53, 70, 247, 15, 171, 66, 128, 218, 71, 210, 226, 175, 85, 102, 77, 81, 242, 178, 195, 123, 204, 248, 116, 143, 227, 37, 23, 151, 141, 55, 215, 84, 112, 92, 172, 136, 190, 217, 138, 14, 113, 147, 47, 28, 206, 144, 252, 241, 73, 162, 48, 91, 224, 52, 58, 65, 157, 212, 72, 3, 222, 185, 193, 166, 231, 234, 165, 101, 
249, 236, 147, 252, 213, 191, 253, 21, 77, 224, 103, 203, 155, 173, 2, 89, 112, 194, 139, 234, 98, 189, 24, 35, 165, 37, 195, 76, 5, 163, 222, 208, 105, 140, 197, 120, 248, 101, 57, 3, 116, 73, 78, 206, 74, 170, 28, 91, 138, 7, 154, 186, 90, 128, 231, 152, 240, 33, 227, 54, 22, 79, 136, 58, 67, 180, 225, 95, 82, 19, 219, 247, 100, 201, 56, 38, 17, 102, 132, 60, 31, 130, 183, 162, 115, 86, 158, 239, 127, 108, 168, 40, 235, 243, 174, 146, 160, 211, 214, 178, 48, 69, 217, 148, 84, 10, 149, 205, 161, 198, 53, 96, 175, 215, 145, 117, 93, 151, 157, 196, 64, 87, 226, 75, 13, 134, 16, 212, 113, 51, 111, 144, 71, 244, 83, 182, 153, 230, 143, 12, 193, 199, 97, 166, 171, 11, 164, 246, 228, 68, 218, 27, 32, 245, 81, 46, 34, 88, 216, 114, 80, 177, 255, 123, 125, 185, 124, 14, 43, 232, 142, 94, 8, 66, 190, 237, 200, 44, 70, 176, 9, 41, 129, 72, 133, 126, 6, 104, 210, 109, 220, 209, 167, 251, 50, 39, 61, 47, 118, 49, 18, 59, 65, 202, 229, 99, 15, 63, 233, 204, 1, 172, 4, 221, 188, 107, 150, 85, 156, 29, 92, 119, 137, 42, 52, 106, 26, 62, 181, 187, 25, 30, 184, 121, 36, 238, 169, 122, 192, 131, 242, 179, 223, 254, 0, 135, 45, 141, 20, 250, 241, 55, 207, 110, 23, 159, 
153, 181, 88, 179, 235, 7, 128, 29, 164, 37, 242, 155, 141, 191, 12, 205, 255, 241, 127, 121, 6, 219, 132, 221, 44, 227, 131, 9, 2, 144, 218, 113, 97, 100, 105, 183, 99, 176, 102, 138, 5, 59, 108, 114, 249, 203, 56, 62, 16, 243, 170, 188, 93, 87, 136, 77, 166, 254, 224, 172, 69, 1, 63, 236, 238, 216, 150, 32, 198, 124, 237, 173, 133, 45, 36, 111, 79, 28, 4, 253, 120, 53, 142, 200, 177, 240, 106, 122, 10, 208, 222, 0, 101, 190, 123, 233, 54, 201, 134, 184, 110, 230, 152, 217, 204, 158, 30, 215, 73, 129, 70, 189, 112, 85, 25, 232, 21, 143, 52, 15, 22, 34, 137, 58, 135, 234, 156, 251, 245, 168, 126, 244, 33, 47, 226, 248, 23, 192, 94, 14, 107, 74, 71, 178, 67, 78, 167, 145, 27, 68, 13, 187, 194, 86, 11, 157, 180, 57, 76, 161, 24, 207, 92, 193, 199, 81, 104, 66, 8, 48, 146, 46, 72, 169, 60, 116, 162, 40, 212, 61, 195, 118, 125, 229, 213, 163, 197, 117, 250, 252, 49, 91, 206, 147, 109, 182, 225, 160, 148, 31, 247, 26, 151, 186, 43, 82, 149, 139, 175, 211, 75, 209, 20, 98, 51, 239, 83, 96, 95, 231, 214, 65, 202, 41, 154, 140, 55, 171, 246, 35, 64, 165, 196, 174, 159, 228, 19, 38, 42, 18, 3, 90, 89, 17, 80, 103, 210, 84, 115, 50, 223, 130, 220, 39, 185, 119, 
130, 206, 255, 207, 242, 227, 122, 205, 193, 80, 99, 10, 252, 164, 128, 144, 146, 235, 42, 189, 106, 76, 135, 140, 31, 197, 249, 57, 239, 48, 7, 168, 69, 142, 248, 151, 63, 253, 167, 89, 6, 114, 214, 229, 234, 52, 220, 123, 88, 129, 40, 102, 224, 93, 94, 111, 231, 222, 137, 75, 101, 11, 243, 172, 103, 237, 208, 165, 200, 178, 45, 188, 177, 109, 157, 126, 154, 190, 124, 72, 187, 54, 181, 26, 201, 185, 104, 100, 120, 198, 143, 183, 1, 221, 131, 79, 118, 32, 47, 161, 245, 236, 215, 65, 160, 66, 35, 191, 68, 4, 85, 92, 116, 210, 108, 147, 141, 3, 39, 87, 84, 145, 223, 61, 113, 174, 78, 250, 19, 202, 44, 175, 64, 18, 33, 115, 77, 228, 9, 209, 132, 55, 51, 0, 83, 24, 97, 180, 121, 53, 43, 213, 29, 67, 119, 204, 195, 184, 163, 149, 139, 134, 176, 13, 186, 166, 70, 251, 95, 27, 158, 90, 218, 5, 127, 196, 50, 219, 199, 226, 179, 241, 217, 240, 62, 23, 211, 169, 171, 58, 96, 192, 8, 37, 30, 49, 73, 117, 74, 98, 16, 254, 28, 153, 182, 133, 247, 212, 246, 107, 81, 105, 170, 155, 216, 38, 156, 244, 125, 138, 173, 194, 82, 22, 150, 59, 41, 46, 232, 17, 71, 12, 60, 36, 34, 152, 230, 136, 159, 21, 15, 20, 112, 110, 2, 86, 56, 225, 91, 238, 148, 233, 203, 25, 162, 14
	);

BEGIN

	-- Instantiate the Unit Under Test (UUT)
	uut: order_perm
	GENERIC MAP(
		DATA_WIDTH => 32,
		M_LOG2 => 8
	)
	PORT MAP(
		clk => clk,
		Dat_in => Dat_in,
		reset => reset,
		datram => datram,
		addr => addr,
		WE => WE,
		Done => Done
	);

	tb : PROCESS
	BEGIN
		wait for clk_T/2;
		clk <= not clk;
	END PROCESS;

	it : process (clk)
	begin
		if (clk = '1' and clk'event) then
			if (done = '0') then
				if (iter = LAST or reset = '1') then
					iter <= 0;
				else
					iter <= iter + 1;
				end if;
			else
				iter <= 0;
			end if;
		end if;
	end process;

	RST:process (clk)
	begin
		if (clk = '1' and clk'event) then
			if (done = '1') then
				reset <= '1';
			else
				reset <= '0';
			end if;
		end if;
	end process;

	--perm_data <= perm_rom(conv_integer(iter));
	perm_data <= perm_rom(iter);
	dat_in <= conv_std_logic_vector(perm_data, 8);

	RA : process (clk)
	begin
		if (clk = '1' and clk'event) then
			if (WE = '1') then
				ram_out(conv_integer(addr)) <= conv_integer(Datram);
			end if;
		end if;
	end process;


END;
